////////////////////////////////////////////////////////////////////-
// Design unit: vm (All In One)
//            :
// File name  : vm.v
//            :
// Description: RTL Design of Vending Machine
//            :
// Limitations: None
//            :
// System     : Verilog
//            :
// Author     : 1. Wan Ahmad Zainie bin Wan Mohamad (ME131135)
//            :    wanahmadzainie@gmail.com
//            : 2. Azfar 'Aizat bin Mohd Isa (ME131032)
//            :    aaizat5@gmail.com
//
// Revision   : Version 0.0 2014-05-30
////////////////////////////////////////////////////////////////////-

module vm(dummy_in, dummy_out);
	input	dummy_in;
	output	dummy_out;

	assign dummy_out = ~dummy_in;
endmodule
