////////////////////////////////////////////////////////////////////-
// Design unit: Control Unit (Module)
//            :
// File name  : cu.v
//            :
// Description: Control Unit of Vending Machine
//            :
// Limitations: None
//            :
// System     : Verilog
//            :
// Author     : Wan Ahmad Zainie bin Wan Mohamad
//            : ME131135
//            : wanahmadzainie@gmail.com
//
// Revision   : Version 0.0 2014-05-30
////////////////////////////////////////////////////////////////////-

module cu(dummy_in, dummy_out);
	input	dummy_in;
	output	dummy_out;

	assign dummy_out = ~dummy_in;
endmodule
